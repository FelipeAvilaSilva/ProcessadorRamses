library verilog;
use verilog.vl_types.all;
entity Ramses_vlg_check_tst is
    port(
        testeValorEnd   : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Ramses_vlg_check_tst;
